--VHDL code of exact multiplier, EM-2 
LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY EM2 IS 
	PORT
	(
		a0 :  IN  STD_LOGIC;
		b0 :  IN  STD_LOGIC;
		a1 :  IN  STD_LOGIC;
		a2 :  IN  STD_LOGIC;
		a3 :  IN  STD_LOGIC;
		a4 :  IN  STD_LOGIC;
		a5 :  IN  STD_LOGIC;
		a6 :  IN  STD_LOGIC;
		a7 :  IN  STD_LOGIC;
		b1 :  IN  STD_LOGIC;
		b2 :  IN  STD_LOGIC;
		b3 :  IN  STD_LOGIC;
		b4 :  IN  STD_LOGIC;
		b5 :  IN  STD_LOGIC;
		b6 :  IN  STD_LOGIC;
		b7 :  IN  STD_LOGIC;
		Low :  IN  STD_LOGIC;
		p0 :  OUT  STD_LOGIC;
		p1 :  OUT  STD_LOGIC;
		p2 :  OUT  STD_LOGIC;
		p3 :  OUT  STD_LOGIC;
		p4 :  OUT  STD_LOGIC;
		p5 :  OUT  STD_LOGIC;
		p6 :  OUT  STD_LOGIC;
		p7 :  OUT  STD_LOGIC;
		p8 :  OUT  STD_LOGIC;
		p9 :  OUT  STD_LOGIC;
		p10 :  OUT  STD_LOGIC;
		p11 :  OUT  STD_LOGIC;
		p12 :  OUT  STD_LOGIC;
		p13 :  OUT  STD_LOGIC;
		p14 :  OUT  STD_LOGIC;
		p15 :  OUT  STD_LOGIC
	);
END EM2;

ARCHITECTURE bdf_type OF EM2 IS 
--component declaration of EFA
COMPONENT fa_opt1
	PORT(bf : IN STD_LOGIC;
		 af : IN STD_LOGIC;
		 c1 : IN STD_LOGIC;
		 sf : OUT STD_LOGIC;
		 cf : OUT STD_LOGIC
	);
END COMPONENT;
--component declaration of IOC
COMPONENT fa_inv1
	PORT(b : IN STD_LOGIC;
		 a : IN STD_LOGIC;
		 ci : IN STD_LOGIC;
		 co : OUT STD_LOGIC;
		 s : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT nands2
	PORT(i1 : IN STD_LOGIC;
		 i2 : IN STD_LOGIC;
		 o1 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT ors2
	PORT(i1 : IN STD_LOGIC;
		 i2 : IN STD_LOGIC;
		 o1 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT ands2
	PORT(i1 : IN STD_LOGIC;
		 i2 : IN STD_LOGIC;
		 o1 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT nots
	PORT(Ai : IN STD_LOGIC;
		 Yi : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT nors2
	PORT(i1 : IN STD_LOGIC;
		 i2 : IN STD_LOGIC;
		 o1 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT nands3
	PORT(i1 : IN STD_LOGIC;
		 i2 : IN STD_LOGIC;
		 i3 : IN STD_LOGIC;
		 o1 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT nands4
	PORT(i1 : IN STD_LOGIC;
		 i2 : IN STD_LOGIC;
		 i3 : IN STD_LOGIC;
		 i4 : IN STD_LOGIC;
		 o1 : OUT STD_LOGIC
	);
END COMPONENT;

--component declaration of IIC
COMPONENT fa_inv
	PORT(b : IN STD_LOGIC;
		 a : IN STD_LOGIC;
		 ci : IN STD_LOGIC;
		 co : OUT STD_LOGIC;
		 s : OUT STD_LOGIC
	);
END COMPONENT;
--component declaration of inverting input half adder
COMPONENT ha_invin1
	PORT(ahc : IN STD_LOGIC;
		 bhc : IN STD_LOGIC;
		 hc : OUT STD_LOGIC;
		 sh : OUT STD_LOGIC
	);
END COMPONENT;
--component declaration of half adder
COMPONENT haxor1
	PORT(bh : IN STD_LOGIC;
		 ah : IN STD_LOGIC;
		 hc : OUT STD_LOGIC;
		 sh : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_354 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_355 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_356 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_357 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_358 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_359 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_360 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_361 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_362 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_363 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_364 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_365 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_366 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_367 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_368 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_369 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_370 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_371 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_372 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_373 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_374 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_375 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_376 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_377 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_378 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_379 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_80 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_380 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_381 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_84 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_382 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_383 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_384 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_385 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_386 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_387 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_388 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_389 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_104 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_390 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_108 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_391 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_112 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_392 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_120 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_393 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_394 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_123 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_124 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_125 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_126 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_127 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_128 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_395 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_396 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_397 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_398 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_399 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_400 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_401 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_145 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_146 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_402 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_403 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_149 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_150 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_151 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_404 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_405 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_406 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_407 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_160 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_161 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_162 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_408 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_409 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_410 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_169 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_411 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_412 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_413 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_177 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_414 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_181 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_415 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_187 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_416 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_417 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_418 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_419 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_420 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_200 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_201 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_202 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_203 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_204 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_206 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_207 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_208 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_209 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_211 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_212 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_213 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_214 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_215 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_216 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_217 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_421 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_422 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_221 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_222 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_223 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_224 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_226 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_227 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_228 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_229 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_230 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_231 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_232 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_234 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_235 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_236 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_237 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_238 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_239 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_243 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_244 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_245 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_246 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_247 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_248 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_249 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_250 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_251 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_256 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_257 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_258 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_260 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_262 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_263 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_264 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_265 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_266 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_267 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_268 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_269 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_270 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_271 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_272 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_273 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_274 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_275 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_276 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_277 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_278 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_279 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_280 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_281 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_282 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_283 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_284 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_285 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_286 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_287 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_288 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_289 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_290 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_291 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_292 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_293 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_294 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_295 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_296 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_297 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_298 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_299 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_300 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_301 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_302 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_303 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_304 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_305 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_306 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_307 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_308 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_309 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_310 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_311 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_312 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_313 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_314 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_315 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_316 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_317 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_318 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_319 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_320 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_321 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_322 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_323 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_324 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_325 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_326 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_327 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_328 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_329 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_330 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_331 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_332 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_333 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_334 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_335 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_336 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_337 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_338 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_339 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_342 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_343 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_346 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_347 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_348 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_349 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_352 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_353 :  STD_LOGIC;


BEGIN 



b2v_inst : fa_opt1
PORT MAP(bf => SYNTHESIZED_WIRE_0,
		 af => SYNTHESIZED_WIRE_1,
		 c1 => SYNTHESIZED_WIRE_2,
		 sf => p4,
		 cf => SYNTHESIZED_WIRE_162);


b2v_inst1 : fa_opt1
PORT MAP(bf => SYNTHESIZED_WIRE_3,
		 af => SYNTHESIZED_WIRE_4,
		 c1 => SYNTHESIZED_WIRE_5,
		 sf => SYNTHESIZED_WIRE_161,
		 cf => SYNTHESIZED_WIRE_208);


b2v_inst10 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_6,
		 a => SYNTHESIZED_WIRE_7,
		 ci => SYNTHESIZED_WIRE_8,
		 co => SYNTHESIZED_WIRE_282,
		 s => SYNTHESIZED_WIRE_277);


b2v_inst11 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_9,
		 a => SYNTHESIZED_WIRE_10,
		 ci => SYNTHESIZED_WIRE_11,
		 co => SYNTHESIZED_WIRE_313,
		 s => SYNTHESIZED_WIRE_280);


b2v_inst12 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_12,
		 a => SYNTHESIZED_WIRE_13,
		 ci => SYNTHESIZED_WIRE_14,
		 co => SYNTHESIZED_WIRE_294,
		 s => SYNTHESIZED_WIRE_289);


b2v_inst121 : nands2
PORT MAP(i1 => b0,
		 i2 => a6,
		 o1 => SYNTHESIZED_WIRE_8);


b2v_inst125 : nands2
PORT MAP(i1 => b4,
		 i2 => a6,
		 o1 => SYNTHESIZED_WIRE_63);


b2v_inst13 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_15,
		 a => SYNTHESIZED_WIRE_16,
		 ci => SYNTHESIZED_WIRE_17,
		 co => SYNTHESIZED_WIRE_297,
		 s => SYNTHESIZED_WIRE_292);


b2v_inst1332 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_354,
		 i2 => SYNTHESIZED_WIRE_355,
		 o1 => SYNTHESIZED_WIRE_357);


b2v_inst1333 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_354,
		 i2 => SYNTHESIZED_WIRE_355,
		 o1 => SYNTHESIZED_WIRE_356);


b2v_inst1334 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_356,
		 i2 => SYNTHESIZED_WIRE_357,
		 o1 => SYNTHESIZED_WIRE_369);


b2v_inst1335 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_358,
		 i2 => SYNTHESIZED_WIRE_356,
		 o1 => SYNTHESIZED_WIRE_26);


b2v_inst1336 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_26,
		 i2 => SYNTHESIZED_WIRE_357,
		 o1 => SYNTHESIZED_WIRE_361);


b2v_inst1337 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_359,
		 i2 => SYNTHESIZED_WIRE_356,
		 o1 => SYNTHESIZED_WIRE_31);


b2v_inst1338 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_360,
		 i2 => SYNTHESIZED_WIRE_31,
		 o1 => SYNTHESIZED_WIRE_362);


b2v_inst1339 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_361,
		 i2 => SYNTHESIZED_WIRE_362,
		 o1 => SYNTHESIZED_WIRE_415);


b2v_inst1340 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_363,
		 i2 => SYNTHESIZED_WIRE_364,
		 o1 => SYNTHESIZED_WIRE_413);


b2v_inst1347 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_365,
		 i2 => SYNTHESIZED_WIRE_366,
		 o1 => SYNTHESIZED_WIRE_367);


b2v_inst1348 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_365,
		 i2 => SYNTHESIZED_WIRE_366,
		 o1 => SYNTHESIZED_WIRE_359);


b2v_inst1349 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_359,
		 i2 => SYNTHESIZED_WIRE_367,
		 o1 => SYNTHESIZED_WIRE_368);


b2v_inst1350 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_366,
		 i2 => SYNTHESIZED_WIRE_365,
		 o1 => SYNTHESIZED_WIRE_358);


b2v_inst1357 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_44,
		 i2 => SYNTHESIZED_WIRE_367,
		 o1 => SYNTHESIZED_WIRE_50);


b2v_inst1363 : nots
PORT MAP(Ai => SYNTHESIZED_WIRE_359,
		 Yi => SYNTHESIZED_WIRE_44);


b2v_inst1376 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_47,
		 i2 => SYNTHESIZED_WIRE_48,
		 o1 => p11);


b2v_inst1379 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_360,
		 i2 => SYNTHESIZED_WIRE_50,
		 o1 => SYNTHESIZED_WIRE_232);


b2v_inst1381 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_51,
		 i2 => SYNTHESIZED_WIRE_52,
		 o1 => p6);


b2v_inst1383 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_53,
		 i2 => SYNTHESIZED_WIRE_54,
		 o1 => p8);


b2v_inst1396 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_360,
		 i2 => SYNTHESIZED_WIRE_368,
		 o1 => SYNTHESIZED_WIRE_52);


b2v_inst1397 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_360,
		 i2 => SYNTHESIZED_WIRE_368,
		 o1 => SYNTHESIZED_WIRE_51);


b2v_inst1399 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_369,
		 i2 => SYNTHESIZED_WIRE_370,
		 o1 => SYNTHESIZED_WIRE_146);


b2v_inst14 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_61,
		 a => SYNTHESIZED_WIRE_62,
		 ci => SYNTHESIZED_WIRE_63,
		 co => SYNTHESIZED_WIRE_300,
		 s => SYNTHESIZED_WIRE_295);


b2v_inst1400 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_369,
		 i2 => SYNTHESIZED_WIRE_370,
		 o1 => SYNTHESIZED_WIRE_145);


b2v_inst1414 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_371,
		 i2 => SYNTHESIZED_WIRE_372,
		 o1 => SYNTHESIZED_WIRE_374);


b2v_inst1415 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_371,
		 i2 => SYNTHESIZED_WIRE_372,
		 o1 => SYNTHESIZED_WIRE_373);


b2v_inst1416 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_373,
		 i2 => SYNTHESIZED_WIRE_374,
		 o1 => SYNTHESIZED_WIRE_395);


b2v_inst1417 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_375,
		 i2 => SYNTHESIZED_WIRE_376,
		 o1 => SYNTHESIZED_WIRE_378);


b2v_inst1418 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_375,
		 i2 => SYNTHESIZED_WIRE_376,
		 o1 => SYNTHESIZED_WIRE_377);


b2v_inst1419 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_377,
		 i2 => SYNTHESIZED_WIRE_378,
		 o1 => SYNTHESIZED_WIRE_396);


b2v_inst1420 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_379,
		 i2 => SYNTHESIZED_WIRE_377,
		 o1 => SYNTHESIZED_WIRE_80);


b2v_inst1421 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_80,
		 i2 => SYNTHESIZED_WIRE_378,
		 o1 => SYNTHESIZED_WIRE_380);


b2v_inst1422 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_380,
		 i2 => SYNTHESIZED_WIRE_381,
		 o1 => SYNTHESIZED_WIRE_84);


b2v_inst1423 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_84,
		 i2 => SYNTHESIZED_WIRE_382,
		 o1 => SYNTHESIZED_WIRE_385);


b2v_inst1424 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_383,
		 i2 => SYNTHESIZED_WIRE_384,
		 o1 => SYNTHESIZED_WIRE_382);


b2v_inst1425 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_383,
		 i2 => SYNTHESIZED_WIRE_384,
		 o1 => SYNTHESIZED_WIRE_381);


b2v_inst1426 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_381,
		 i2 => SYNTHESIZED_WIRE_382,
		 o1 => SYNTHESIZED_WIRE_399);


b2v_inst1427 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_385,
		 i2 => SYNTHESIZED_WIRE_386,
		 o1 => SYNTHESIZED_WIRE_94);


b2v_inst1428 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_94,
		 i2 => SYNTHESIZED_WIRE_387,
		 o1 => SYNTHESIZED_WIRE_348);


b2v_inst1429 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_388,
		 i2 => SYNTHESIZED_WIRE_389,
		 o1 => SYNTHESIZED_WIRE_387);


b2v_inst1430 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_388,
		 i2 => SYNTHESIZED_WIRE_389,
		 o1 => SYNTHESIZED_WIRE_386);


b2v_inst1431 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_386,
		 i2 => SYNTHESIZED_WIRE_387,
		 o1 => SYNTHESIZED_WIRE_401);


b2v_inst1436 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_372,
		 i2 => SYNTHESIZED_WIRE_371,
		 o1 => SYNTHESIZED_WIRE_379);


b2v_inst1449 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_104,
		 i2 => SYNTHESIZED_WIRE_374,
		 o1 => SYNTHESIZED_WIRE_390);


b2v_inst1450 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_390,
		 i2 => SYNTHESIZED_WIRE_377,
		 o1 => SYNTHESIZED_WIRE_108);


b2v_inst1451 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_108,
		 i2 => SYNTHESIZED_WIRE_378,
		 o1 => SYNTHESIZED_WIRE_391);


b2v_inst1452 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_391,
		 i2 => SYNTHESIZED_WIRE_381,
		 o1 => SYNTHESIZED_WIRE_112);


b2v_inst1453 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_112,
		 i2 => SYNTHESIZED_WIRE_382,
		 o1 => SYNTHESIZED_WIRE_120);


b2v_inst1455 : nots
PORT MAP(Ai => SYNTHESIZED_WIRE_373,
		 Yi => SYNTHESIZED_WIRE_104);


b2v_inst1470 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_392,
		 i2 => SYNTHESIZED_WIRE_390,
		 o1 => SYNTHESIZED_WIRE_209);


b2v_inst1472 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_392,
		 i2 => SYNTHESIZED_WIRE_391,
		 o1 => SYNTHESIZED_WIRE_217);


b2v_inst1474 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_392,
		 i2 => SYNTHESIZED_WIRE_120,
		 o1 => SYNTHESIZED_WIRE_224);


b2v_inst1475 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_393,
		 i2 => SYNTHESIZED_WIRE_394,
		 o1 => SYNTHESIZED_WIRE_352);


b2v_inst1477 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_123,
		 i2 => SYNTHESIZED_WIRE_124,
		 o1 => p14);


b2v_inst1479 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_125,
		 i2 => SYNTHESIZED_WIRE_126,
		 o1 => p13);


b2v_inst1481 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_127,
		 i2 => SYNTHESIZED_WIRE_128,
		 o1 => p12);


b2v_inst1483 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_392,
		 i2 => SYNTHESIZED_WIRE_395,
		 o1 => SYNTHESIZED_WIRE_48);


b2v_inst1484 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_392,
		 i2 => SYNTHESIZED_WIRE_395,
		 o1 => SYNTHESIZED_WIRE_47);


b2v_inst1486 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_396,
		 i2 => SYNTHESIZED_WIRE_397,
		 o1 => SYNTHESIZED_WIRE_128);


b2v_inst1487 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_396,
		 i2 => SYNTHESIZED_WIRE_397,
		 o1 => SYNTHESIZED_WIRE_127);


b2v_inst1489 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_398,
		 i2 => SYNTHESIZED_WIRE_399,
		 o1 => SYNTHESIZED_WIRE_126);


b2v_inst149 : nands2
PORT MAP(i1 => b1,
		 i2 => a5,
		 o1 => SYNTHESIZED_WIRE_7);


b2v_inst1490 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_398,
		 i2 => SYNTHESIZED_WIRE_399,
		 o1 => SYNTHESIZED_WIRE_125);


b2v_inst1492 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_400,
		 i2 => SYNTHESIZED_WIRE_401,
		 o1 => SYNTHESIZED_WIRE_124);


b2v_inst1493 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_400,
		 i2 => SYNTHESIZED_WIRE_401,
		 o1 => SYNTHESIZED_WIRE_123);


b2v_inst1494 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_145,
		 i2 => SYNTHESIZED_WIRE_146,
		 o1 => p7);


b2v_inst1497 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_402,
		 i2 => SYNTHESIZED_WIRE_403,
		 o1 => SYNTHESIZED_WIRE_405);


b2v_inst15 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_149,
		 a => SYNTHESIZED_WIRE_150,
		 ci => SYNTHESIZED_WIRE_151,
		 co => SYNTHESIZED_WIRE_320,
		 s => SYNTHESIZED_WIRE_298);


b2v_inst150 : nands2
PORT MAP(i1 => b1,
		 i2 => a6,
		 o1 => SYNTHESIZED_WIRE_10);


b2v_inst1500 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_402,
		 i2 => SYNTHESIZED_WIRE_403,
		 o1 => SYNTHESIZED_WIRE_404);


b2v_inst1503 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_404,
		 i2 => SYNTHESIZED_WIRE_405,
		 o1 => SYNTHESIZED_WIRE_416);


b2v_inst1504 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_403,
		 i2 => SYNTHESIZED_WIRE_402,
		 o1 => SYNTHESIZED_WIRE_410);


b2v_inst1506 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_406,
		 i2 => SYNTHESIZED_WIRE_407,
		 o1 => SYNTHESIZED_WIRE_409);


b2v_inst151 : nands2
PORT MAP(i1 => b2,
		 i2 => a5,
		 o1 => SYNTHESIZED_WIRE_9);


b2v_inst152 : nands2
PORT MAP(i1 => b2,
		 i2 => a6,
		 o1 => SYNTHESIZED_WIRE_256);


b2v_inst153 : nands2
PORT MAP(i1 => b0,
		 i2 => a5,
		 o1 => SYNTHESIZED_WIRE_276);


b2v_inst154 : nands2
PORT MAP(i1 => b0,
		 i2 => a4,
		 o1 => SYNTHESIZED_WIRE_264);


b2v_inst155 : nands2
PORT MAP(i1 => b0,
		 i2 => a3,
		 o1 => SYNTHESIZED_WIRE_248);


b2v_inst156 : nands2
PORT MAP(i1 => b0,
		 i2 => a2,
		 o1 => SYNTHESIZED_WIRE_216);


b2v_inst157 : nands2
PORT MAP(i1 => b0,
		 i2 => a1,
		 o1 => SYNTHESIZED_WIRE_302);


b2v_inst158 : nands2
PORT MAP(i1 => b1,
		 i2 => a0,
		 o1 => SYNTHESIZED_WIRE_301);


b2v_inst159 : nands2
PORT MAP(i1 => b2,
		 i2 => a0,
		 o1 => SYNTHESIZED_WIRE_214);


b2v_inst16 : fa_opt1
PORT MAP(bf => SYNTHESIZED_WIRE_160,
		 af => SYNTHESIZED_WIRE_161,
		 c1 => SYNTHESIZED_WIRE_162,
		 sf => p5,
		 cf => SYNTHESIZED_WIRE_360);


b2v_inst160 : nands2
PORT MAP(i1 => b1,
		 i2 => a1,
		 o1 => SYNTHESIZED_WIRE_215);


b2v_inst161 : nands2
PORT MAP(i1 => b1,
		 i2 => a2,
		 o1 => SYNTHESIZED_WIRE_247);


b2v_inst162 : nands2
PORT MAP(i1 => b1,
		 i2 => a3,
		 o1 => SYNTHESIZED_WIRE_263);


b2v_inst163 : nands2
PORT MAP(i1 => b1,
		 i2 => a4,
		 o1 => SYNTHESIZED_WIRE_275);


b2v_inst164 : nands2
PORT MAP(i1 => b2,
		 i2 => a3,
		 o1 => SYNTHESIZED_WIRE_274);


b2v_inst165 : nands2
PORT MAP(i1 => b2,
		 i2 => a4,
		 o1 => SYNTHESIZED_WIRE_6);


b2v_inst166 : nands2
PORT MAP(i1 => b2,
		 i2 => a2,
		 o1 => SYNTHESIZED_WIRE_262);


b2v_inst1667 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_406,
		 i2 => SYNTHESIZED_WIRE_407,
		 o1 => SYNTHESIZED_WIRE_408);


b2v_inst1668 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_408,
		 i2 => SYNTHESIZED_WIRE_409,
		 o1 => SYNTHESIZED_WIRE_417);


b2v_inst1669 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_410,
		 i2 => SYNTHESIZED_WIRE_408,
		 o1 => SYNTHESIZED_WIRE_169);


b2v_inst167 : nands2
PORT MAP(i1 => b2,
		 i2 => a1,
		 o1 => SYNTHESIZED_WIRE_246);


b2v_inst1670 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_169,
		 i2 => SYNTHESIZED_WIRE_409,
		 o1 => SYNTHESIZED_WIRE_411);


b2v_inst1671 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_411,
		 i2 => SYNTHESIZED_WIRE_412,
		 o1 => SYNTHESIZED_WIRE_204);


b2v_inst1672 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_363,
		 i2 => SYNTHESIZED_WIRE_364,
		 o1 => SYNTHESIZED_WIRE_412);


b2v_inst1673 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_412,
		 i2 => SYNTHESIZED_WIRE_413,
		 o1 => SYNTHESIZED_WIRE_420);


b2v_inst1674 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_177,
		 i2 => SYNTHESIZED_WIRE_405,
		 o1 => SYNTHESIZED_WIRE_414);


b2v_inst1675 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_414,
		 i2 => SYNTHESIZED_WIRE_408,
		 o1 => SYNTHESIZED_WIRE_181);


b2v_inst1676 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_181,
		 i2 => SYNTHESIZED_WIRE_409,
		 o1 => SYNTHESIZED_WIRE_187);


b2v_inst1679 : nots
PORT MAP(Ai => SYNTHESIZED_WIRE_404,
		 Yi => SYNTHESIZED_WIRE_177);


b2v_inst168 : nands2
PORT MAP(i1 => b5,
		 i2 => a5,
		 o1 => SYNTHESIZED_WIRE_62);


b2v_inst1680 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_415,
		 i2 => SYNTHESIZED_WIRE_414,
		 o1 => SYNTHESIZED_WIRE_258);


b2v_inst1681 : ands2
PORT MAP(i1 => SYNTHESIZED_WIRE_415,
		 i2 => SYNTHESIZED_WIRE_187,
		 o1 => SYNTHESIZED_WIRE_260);


b2v_inst1682 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_415,
		 i2 => SYNTHESIZED_WIRE_416,
		 o1 => SYNTHESIZED_WIRE_54);


b2v_inst1683 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_415,
		 i2 => SYNTHESIZED_WIRE_416,
		 o1 => SYNTHESIZED_WIRE_53);


b2v_inst1684 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_417,
		 i2 => SYNTHESIZED_WIRE_418,
		 o1 => SYNTHESIZED_WIRE_203);


b2v_inst1685 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_417,
		 i2 => SYNTHESIZED_WIRE_418,
		 o1 => SYNTHESIZED_WIRE_202);


b2v_inst1686 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_419,
		 i2 => SYNTHESIZED_WIRE_420,
		 o1 => SYNTHESIZED_WIRE_201);


b2v_inst1687 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_419,
		 i2 => SYNTHESIZED_WIRE_420,
		 o1 => SYNTHESIZED_WIRE_200);


b2v_inst1688 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_200,
		 i2 => SYNTHESIZED_WIRE_201,
		 o1 => p10);


b2v_inst1689 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_202,
		 i2 => SYNTHESIZED_WIRE_203,
		 o1 => p9);


b2v_inst169 : nands2
PORT MAP(i1 => b5,
		 i2 => a6,
		 o1 => SYNTHESIZED_WIRE_150);


b2v_inst1690 : nands2
PORT MAP(i1 => SYNTHESIZED_WIRE_204,
		 i2 => SYNTHESIZED_WIRE_413,
		 o1 => SYNTHESIZED_WIRE_421);


b2v_inst17 : fa_opt1
PORT MAP(bf => SYNTHESIZED_WIRE_206,
		 af => SYNTHESIZED_WIRE_207,
		 c1 => SYNTHESIZED_WIRE_208,
		 sf => SYNTHESIZED_WIRE_365,
		 cf => SYNTHESIZED_WIRE_354);


b2v_inst170 : nands2
PORT MAP(i1 => b6,
		 i2 => a5,
		 o1 => SYNTHESIZED_WIRE_149);


b2v_inst171 : nands2
PORT MAP(i1 => b6,
		 i2 => a6,
		 o1 => SYNTHESIZED_WIRE_315);


b2v_inst172 : nands2
PORT MAP(i1 => b4,
		 i2 => a5,
		 o1 => SYNTHESIZED_WIRE_17);


b2v_inst173 : nands2
PORT MAP(i1 => b4,
		 i2 => a4,
		 o1 => SYNTHESIZED_WIRE_14);


b2v_inst174 : nands2
PORT MAP(i1 => b4,
		 i2 => a3,
		 o1 => SYNTHESIZED_WIRE_339);


b2v_inst175 : nands2
PORT MAP(i1 => b4,
		 i2 => a2,
		 o1 => SYNTHESIZED_WIRE_305);


b2v_inst176 : nands2
PORT MAP(i1 => b4,
		 i2 => a1,
		 o1 => SYNTHESIZED_WIRE_307);


b2v_inst177 : nands2
PORT MAP(i1 => b5,
		 i2 => a0,
		 o1 => SYNTHESIZED_WIRE_306);


b2v_inst178 : nands2
PORT MAP(i1 => b6,
		 i2 => a0,
		 o1 => SYNTHESIZED_WIRE_303);


b2v_inst179 : nands2
PORT MAP(i1 => b5,
		 i2 => a1,
		 o1 => SYNTHESIZED_WIRE_304);


b2v_inst18 : nors2
PORT MAP(i1 => SYNTHESIZED_WIRE_209,
		 i2 => SYNTHESIZED_WIRE_379,
		 o1 => SYNTHESIZED_WIRE_397);


b2v_inst180 : nands2
PORT MAP(i1 => b5,
		 i2 => a2,
		 o1 => SYNTHESIZED_WIRE_338);


b2v_inst181 : nands2
PORT MAP(i1 => b5,
		 i2 => a3,
		 o1 => SYNTHESIZED_WIRE_13);


b2v_inst182 : nands2
PORT MAP(i1 => b5,
		 i2 => a4,
		 o1 => SYNTHESIZED_WIRE_16);


b2v_inst183 : nands2
PORT MAP(i1 => b6,
		 i2 => a3,
		 o1 => SYNTHESIZED_WIRE_15);


b2v_inst184 : nands2
PORT MAP(i1 => b6,
		 i2 => a4,
		 o1 => SYNTHESIZED_WIRE_61);


b2v_inst185 : nands2
PORT MAP(i1 => b6,
		 i2 => a2,
		 o1 => SYNTHESIZED_WIRE_12);


b2v_inst186 : nands2
PORT MAP(i1 => b6,
		 i2 => a1,
		 o1 => SYNTHESIZED_WIRE_337);


b2v_inst189 : nands2
PORT MAP(i1 => b3,
		 i2 => a0,
		 o1 => SYNTHESIZED_WIRE_266);


b2v_inst19 : fa_opt1
PORT MAP(bf => SYNTHESIZED_WIRE_211,
		 af => SYNTHESIZED_WIRE_212,
		 c1 => SYNTHESIZED_WIRE_213,
		 sf => SYNTHESIZED_WIRE_355,
		 cf => SYNTHESIZED_WIRE_402);


b2v_inst190 : nands2
PORT MAP(i1 => b3,
		 i2 => a1,
		 o1 => SYNTHESIZED_WIRE_269);


b2v_inst191 : nands2
PORT MAP(i1 => b3,
		 i2 => a3,
		 o1 => SYNTHESIZED_WIRE_278);


b2v_inst192 : nands2
PORT MAP(i1 => b3,
		 i2 => a2,
		 o1 => SYNTHESIZED_WIRE_272);


b2v_inst194 : nands2
PORT MAP(i1 => b3,
		 i2 => a4,
		 o1 => SYNTHESIZED_WIRE_281);


b2v_inst195 : nands2
PORT MAP(i1 => b3,
		 i2 => a5,
		 o1 => SYNTHESIZED_WIRE_311);


b2v_inst196 : nands2
PORT MAP(i1 => b3,
		 i2 => a6,
		 o1 => SYNTHESIZED_WIRE_283);


b2v_inst197 : nands2
PORT MAP(i1 => b3,
		 i2 => a7,
		 o1 => SYNTHESIZED_WIRE_243);


b2v_inst2 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_214,
		 a => SYNTHESIZED_WIRE_215,
		 ci => SYNTHESIZED_WIRE_216,
		 co => SYNTHESIZED_WIRE_267,
		 s => SYNTHESIZED_WIRE_314);


b2v_inst20 : nors2
PORT MAP(i1 => SYNTHESIZED_WIRE_217,
		 i2 => SYNTHESIZED_WIRE_380,
		 o1 => SYNTHESIZED_WIRE_398);


b2v_inst2057 : ors2
PORT MAP(i1 => SYNTHESIZED_WIRE_421,
		 i2 => SYNTHESIZED_WIRE_422,
		 o1 => SYNTHESIZED_WIRE_392);


b2v_inst21 : fa_opt1
PORT MAP(bf => SYNTHESIZED_WIRE_221,
		 af => SYNTHESIZED_WIRE_222,
		 c1 => SYNTHESIZED_WIRE_223,
		 sf => SYNTHESIZED_WIRE_403,
		 cf => SYNTHESIZED_WIRE_406);


b2v_inst22 : nors2
PORT MAP(i1 => SYNTHESIZED_WIRE_224,
		 i2 => SYNTHESIZED_WIRE_385,
		 o1 => SYNTHESIZED_WIRE_400);


b2v_inst23 : fa_opt1
PORT MAP(bf => SYNTHESIZED_WIRE_226,
		 af => SYNTHESIZED_WIRE_227,
		 c1 => SYNTHESIZED_WIRE_228,
		 sf => SYNTHESIZED_WIRE_221,
		 cf => SYNTHESIZED_WIRE_230);


b2v_inst24 : fa_opt1
PORT MAP(bf => SYNTHESIZED_WIRE_229,
		 af => SYNTHESIZED_WIRE_230,
		 c1 => SYNTHESIZED_WIRE_231,
		 sf => SYNTHESIZED_WIRE_407,
		 cf => SYNTHESIZED_WIRE_364);


b2v_inst25 : nors2
PORT MAP(i1 => SYNTHESIZED_WIRE_232,
		 i2 => SYNTHESIZED_WIRE_358,
		 o1 => SYNTHESIZED_WIRE_370);


b2v_inst26 : fa_opt1
PORT MAP(bf => SYNTHESIZED_WIRE_234,
		 af => SYNTHESIZED_WIRE_235,
		 c1 => SYNTHESIZED_WIRE_236,
		 sf => SYNTHESIZED_WIRE_229,
		 cf => SYNTHESIZED_WIRE_238);


b2v_inst27 : fa_opt1
PORT MAP(bf => SYNTHESIZED_WIRE_237,
		 af => SYNTHESIZED_WIRE_238,
		 c1 => SYNTHESIZED_WIRE_239,
		 sf => SYNTHESIZED_WIRE_363,
		 cf => SYNTHESIZED_WIRE_371);


b2v_inst28 : nands3
PORT MAP(i1 => SYNTHESIZED_WIRE_404,
		 i2 => SYNTHESIZED_WIRE_408,
		 i3 => SYNTHESIZED_WIRE_412,
		 o1 => SYNTHESIZED_WIRE_343);


b2v_inst29 : fa_opt1
PORT MAP(bf => SYNTHESIZED_WIRE_243,
		 af => SYNTHESIZED_WIRE_244,
		 c1 => SYNTHESIZED_WIRE_245,
		 sf => SYNTHESIZED_WIRE_237,
		 cf => SYNTHESIZED_WIRE_250);


b2v_inst3 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_246,
		 a => SYNTHESIZED_WIRE_247,
		 ci => SYNTHESIZED_WIRE_248,
		 co => SYNTHESIZED_WIRE_270,
		 s => SYNTHESIZED_WIRE_265);


b2v_inst30 : fa_opt1
PORT MAP(bf => SYNTHESIZED_WIRE_249,
		 af => SYNTHESIZED_WIRE_250,
		 c1 => SYNTHESIZED_WIRE_251,
		 sf => SYNTHESIZED_WIRE_372,
		 cf => SYNTHESIZED_WIRE_375);


b2v_inst31 : nands4
PORT MAP(i1 => SYNTHESIZED_WIRE_373,
		 i2 => SYNTHESIZED_WIRE_377,
		 i3 => SYNTHESIZED_WIRE_381,
		 i4 => SYNTHESIZED_WIRE_386,
		 o1 => SYNTHESIZED_WIRE_347);


b2v_inst32 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_256,
		 a => SYNTHESIZED_WIRE_257,
		 ci => Low,
		 co => SYNTHESIZED_WIRE_285,
		 s => SYNTHESIZED_WIRE_312);


b2v_inst36 : nors2
PORT MAP(i1 => SYNTHESIZED_WIRE_258,
		 i2 => SYNTHESIZED_WIRE_410,
		 o1 => SYNTHESIZED_WIRE_418);


b2v_inst37 : nors2
PORT MAP(i1 => SYNTHESIZED_WIRE_260,
		 i2 => SYNTHESIZED_WIRE_411,
		 o1 => SYNTHESIZED_WIRE_419);


b2v_inst4 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_262,
		 a => SYNTHESIZED_WIRE_263,
		 ci => SYNTHESIZED_WIRE_264,
		 co => SYNTHESIZED_WIRE_273,
		 s => SYNTHESIZED_WIRE_268);


b2v_inst47 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_265,
		 a => SYNTHESIZED_WIRE_266,
		 ci => SYNTHESIZED_WIRE_267,
		 co => SYNTHESIZED_WIRE_327,
		 s => SYNTHESIZED_WIRE_326);


b2v_inst48 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_268,
		 a => SYNTHESIZED_WIRE_269,
		 ci => SYNTHESIZED_WIRE_270,
		 co => SYNTHESIZED_WIRE_4,
		 s => SYNTHESIZED_WIRE_328);


b2v_inst49 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_271,
		 a => SYNTHESIZED_WIRE_272,
		 ci => SYNTHESIZED_WIRE_273,
		 co => SYNTHESIZED_WIRE_207,
		 s => SYNTHESIZED_WIRE_3);


b2v_inst5 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_274,
		 a => SYNTHESIZED_WIRE_275,
		 ci => SYNTHESIZED_WIRE_276,
		 co => SYNTHESIZED_WIRE_279,
		 s => SYNTHESIZED_WIRE_271);


b2v_inst50 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_277,
		 a => SYNTHESIZED_WIRE_278,
		 ci => SYNTHESIZED_WIRE_279,
		 co => SYNTHESIZED_WIRE_329,
		 s => SYNTHESIZED_WIRE_206);


b2v_inst51 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_280,
		 a => SYNTHESIZED_WIRE_281,
		 ci => SYNTHESIZED_WIRE_282,
		 co => SYNTHESIZED_WIRE_227,
		 s => SYNTHESIZED_WIRE_330);


b2v_inst52 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_283,
		 a => SYNTHESIZED_WIRE_284,
		 ci => SYNTHESIZED_WIRE_285,
		 co => SYNTHESIZED_WIRE_244,
		 s => SYNTHESIZED_WIRE_234);


b2v_inst54 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_286,
		 a => SYNTHESIZED_WIRE_287,
		 ci => SYNTHESIZED_WIRE_288,
		 co => SYNTHESIZED_WIRE_228,
		 s => SYNTHESIZED_WIRE_213);


b2v_inst55 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_289,
		 a => SYNTHESIZED_WIRE_290,
		 ci => SYNTHESIZED_WIRE_291,
		 co => SYNTHESIZED_WIRE_236,
		 s => SYNTHESIZED_WIRE_223);


b2v_inst56 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_292,
		 a => SYNTHESIZED_WIRE_293,
		 ci => SYNTHESIZED_WIRE_294,
		 co => SYNTHESIZED_WIRE_245,
		 s => SYNTHESIZED_WIRE_231);


b2v_inst57 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_295,
		 a => SYNTHESIZED_WIRE_296,
		 ci => SYNTHESIZED_WIRE_297,
		 co => SYNTHESIZED_WIRE_249,
		 s => SYNTHESIZED_WIRE_239);


b2v_inst58 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_298,
		 a => SYNTHESIZED_WIRE_299,
		 ci => SYNTHESIZED_WIRE_300,
		 co => SYNTHESIZED_WIRE_332,
		 s => SYNTHESIZED_WIRE_251);


b2v_inst59 : ha_invin1
PORT MAP(ahc => SYNTHESIZED_WIRE_301,
		 bhc => SYNTHESIZED_WIRE_302,
		 hc => SYNTHESIZED_WIRE_318,
		 sh => p1);


b2v_inst6 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_303,
		 a => SYNTHESIZED_WIRE_304,
		 ci => SYNTHESIZED_WIRE_305,
		 co => SYNTHESIZED_WIRE_288,
		 s => SYNTHESIZED_WIRE_322);


b2v_inst60 : ha_invin1
PORT MAP(ahc => SYNTHESIZED_WIRE_306,
		 bhc => SYNTHESIZED_WIRE_307,
		 hc => SYNTHESIZED_WIRE_323,
		 sh => SYNTHESIZED_WIRE_160);


b2v_inst61 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_308,
		 a => SYNTHESIZED_WIRE_309,
		 ci => SYNTHESIZED_WIRE_310,
		 co => SYNTHESIZED_WIRE_336,
		 s => SYNTHESIZED_WIRE_333);


b2v_inst62 : ands2
PORT MAP(i1 => b7,
		 i2 => a7,
		 o1 => SYNTHESIZED_WIRE_335);


b2v_inst63 : ands2
PORT MAP(i1 => b0,
		 i2 => a7,
		 o1 => SYNTHESIZED_WIRE_11);


b2v_inst64 : ands2
PORT MAP(i1 => b1,
		 i2 => a7,
		 o1 => SYNTHESIZED_WIRE_257);


b2v_inst65 : ands2
PORT MAP(i1 => b2,
		 i2 => a7,
		 o1 => SYNTHESIZED_WIRE_284);


b2v_inst66 : ands2
PORT MAP(i1 => b4,
		 i2 => a7,
		 o1 => SYNTHESIZED_WIRE_151);


b2v_inst67 : ands2
PORT MAP(i1 => b5,
		 i2 => a7,
		 o1 => SYNTHESIZED_WIRE_316);


b2v_inst68 : ands2
PORT MAP(i1 => b6,
		 i2 => a7,
		 o1 => SYNTHESIZED_WIRE_309);


b2v_inst69 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_311,
		 a => SYNTHESIZED_WIRE_312,
		 ci => SYNTHESIZED_WIRE_313,
		 co => SYNTHESIZED_WIRE_235,
		 s => SYNTHESIZED_WIRE_226);


b2v_inst7 : ands2
PORT MAP(i1 => b0,
		 i2 => a0,
		 o1 => p0);


b2v_inst71 : nots
PORT MAP(Ai => SYNTHESIZED_WIRE_314,
		 Yi => SYNTHESIZED_WIRE_319);


b2v_inst72 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_315,
		 a => SYNTHESIZED_WIRE_316,
		 ci => SYNTHESIZED_WIRE_317,
		 co => SYNTHESIZED_WIRE_310,
		 s => SYNTHESIZED_WIRE_321);


b2v_inst73 : haxor1
PORT MAP(bh => SYNTHESIZED_WIRE_318,
		 ah => SYNTHESIZED_WIRE_319,
		 hc => SYNTHESIZED_WIRE_325,
		 sh => p2);


b2v_inst74 : ha_invin1
PORT MAP(ahc => SYNTHESIZED_WIRE_320,
		 bhc => SYNTHESIZED_WIRE_321,
		 hc => SYNTHESIZED_WIRE_334,
		 sh => SYNTHESIZED_WIRE_331);


b2v_inst75 : nots
PORT MAP(Ai => SYNTHESIZED_WIRE_322,
		 Yi => SYNTHESIZED_WIRE_324);


b2v_inst76 : haxor1
PORT MAP(bh => SYNTHESIZED_WIRE_323,
		 ah => SYNTHESIZED_WIRE_324,
		 hc => SYNTHESIZED_WIRE_212,
		 sh => SYNTHESIZED_WIRE_366);


b2v_inst77 : haxor1
PORT MAP(bh => SYNTHESIZED_WIRE_325,
		 ah => SYNTHESIZED_WIRE_326,
		 hc => SYNTHESIZED_WIRE_2,
		 sh => p3);


b2v_inst78 : haxor1
PORT MAP(bh => SYNTHESIZED_WIRE_327,
		 ah => SYNTHESIZED_WIRE_328,
		 hc => SYNTHESIZED_WIRE_5,
		 sh => SYNTHESIZED_WIRE_0);


b2v_inst79 : haxor1
PORT MAP(bh => SYNTHESIZED_WIRE_329,
		 ah => SYNTHESIZED_WIRE_330,
		 hc => SYNTHESIZED_WIRE_222,
		 sh => SYNTHESIZED_WIRE_211);


b2v_inst8 : ands2
PORT MAP(i1 => b4,
		 i2 => a0,
		 o1 => SYNTHESIZED_WIRE_1);


b2v_inst80 : haxor1
PORT MAP(bh => SYNTHESIZED_WIRE_331,
		 ah => SYNTHESIZED_WIRE_332,
		 hc => SYNTHESIZED_WIRE_384,
		 sh => SYNTHESIZED_WIRE_376);


b2v_inst81 : haxor1
PORT MAP(bh => SYNTHESIZED_WIRE_333,
		 ah => SYNTHESIZED_WIRE_334,
		 hc => SYNTHESIZED_WIRE_389,
		 sh => SYNTHESIZED_WIRE_383);


b2v_inst82 : haxor1
PORT MAP(bh => SYNTHESIZED_WIRE_335,
		 ah => SYNTHESIZED_WIRE_336,
		 hc => SYNTHESIZED_WIRE_394,
		 sh => SYNTHESIZED_WIRE_388);


b2v_inst83 : ands2
PORT MAP(i1 => b7,
		 i2 => a6,
		 o1 => SYNTHESIZED_WIRE_308);


b2v_inst84 : ands2
PORT MAP(i1 => b7,
		 i2 => a5,
		 o1 => SYNTHESIZED_WIRE_317);


b2v_inst85 : ands2
PORT MAP(i1 => b7,
		 i2 => a4,
		 o1 => SYNTHESIZED_WIRE_299);


b2v_inst86 : ands2
PORT MAP(i1 => b7,
		 i2 => a3,
		 o1 => SYNTHESIZED_WIRE_296);


b2v_inst87 : ands2
PORT MAP(i1 => b7,
		 i2 => a2,
		 o1 => SYNTHESIZED_WIRE_293);


b2v_inst88 : ands2
PORT MAP(i1 => b7,
		 i2 => a1,
		 o1 => SYNTHESIZED_WIRE_290);


b2v_inst89 : ands2
PORT MAP(i1 => b7,
		 i2 => a0,
		 o1 => SYNTHESIZED_WIRE_287);


b2v_inst9 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_337,
		 a => SYNTHESIZED_WIRE_338,
		 ci => SYNTHESIZED_WIRE_339,
		 co => SYNTHESIZED_WIRE_291,
		 s => SYNTHESIZED_WIRE_286);


b2v_inst90 : nors2
PORT MAP(i1 => SYNTHESIZED_WIRE_361,
		 i2 => SYNTHESIZED_WIRE_362,
		 o1 => SYNTHESIZED_WIRE_342);


b2v_inst91 : nors2
PORT MAP(i1 => SYNTHESIZED_WIRE_342,
		 i2 => SYNTHESIZED_WIRE_343,
		 o1 => SYNTHESIZED_WIRE_422);


b2v_inst92 : nors2
PORT MAP(i1 => SYNTHESIZED_WIRE_421,
		 i2 => SYNTHESIZED_WIRE_422,
		 o1 => SYNTHESIZED_WIRE_346);


b2v_inst93 : nors2
PORT MAP(i1 => SYNTHESIZED_WIRE_346,
		 i2 => SYNTHESIZED_WIRE_347,
		 o1 => SYNTHESIZED_WIRE_349);


b2v_inst94 : nors2
PORT MAP(i1 => SYNTHESIZED_WIRE_348,
		 i2 => SYNTHESIZED_WIRE_349,
		 o1 => SYNTHESIZED_WIRE_393);


b2v_inst95 : nors2
PORT MAP(i1 => SYNTHESIZED_WIRE_394,
		 i2 => SYNTHESIZED_WIRE_393,
		 o1 => SYNTHESIZED_WIRE_353);


b2v_inst96 : nors2
PORT MAP(i1 => SYNTHESIZED_WIRE_352,
		 i2 => SYNTHESIZED_WIRE_353,
		 o1 => p15);


END bdf_type;
