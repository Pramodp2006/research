--VHDL code for the approximate multiplier, APM-8
LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY APM8 IS 
	PORT
	(
		a0 :  IN  STD_LOGIC;
		b0 :  IN  STD_LOGIC;
		a1 :  IN  STD_LOGIC;
		a2 :  IN  STD_LOGIC;
		a3 :  IN  STD_LOGIC;
		a4 :  IN  STD_LOGIC;
		a5 :  IN  STD_LOGIC;
		a6 :  IN  STD_LOGIC;
		a7 :  IN  STD_LOGIC;
		b1 :  IN  STD_LOGIC;
		b2 :  IN  STD_LOGIC;
		b3 :  IN  STD_LOGIC;
		b4 :  IN  STD_LOGIC;
		b5 :  IN  STD_LOGIC;
		b6 :  IN  STD_LOGIC;
		b7 :  IN  STD_LOGIC;
		Low :  IN  STD_LOGIC;
		p0 :  OUT  STD_LOGIC;
		p1 :  OUT  STD_LOGIC;
		p2 :  OUT  STD_LOGIC;
		p3 :  OUT  STD_LOGIC;
		p4 :  OUT  STD_LOGIC;
		p5 :  OUT  STD_LOGIC;
		p6 :  OUT  STD_LOGIC;
		p7 :  OUT  STD_LOGIC;
		p8 :  OUT  STD_LOGIC;
		p9 :  OUT  STD_LOGIC;
		p10 :  OUT  STD_LOGIC;
		p11 :  OUT  STD_LOGIC;
		p12 :  OUT  STD_LOGIC;
		p13 :  OUT  STD_LOGIC;
		p14 :  OUT  STD_LOGIC;
		p15 :  OUT  STD_LOGIC
	);
END APM8;

ARCHITECTURE bdf_type OF APM8 IS 
--Component declaration of AOFA-1
COMPONENT fa_inv1app
	PORT(b : IN STD_LOGIC;
		 a : IN STD_LOGIC;
		 ci : IN STD_LOGIC;
		 s : OUT STD_LOGIC;
		 co : OUT STD_LOGIC
	);
END COMPONENT;
--Component declaration of IOC
COMPONENT fa_inv1
	PORT(b : IN STD_LOGIC;
		 a : IN STD_LOGIC;
		 ci : IN STD_LOGIC;
		 co : OUT STD_LOGIC;
		 s : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT nands2
	PORT(i1 : IN STD_LOGIC;
		 i2 : IN STD_LOGIC;
		 o1 : OUT STD_LOGIC
	);
END COMPONENT;
--Component declaration of AIFA-2
COMPONENT fainvimpapp
	PORT(b : IN STD_LOGIC;
		 a : IN STD_LOGIC;
		 ci : IN STD_LOGIC;
		 co : OUT STD_LOGIC;
		 s : OUT STD_LOGIC
	);
END COMPONENT;
--Component declaration of AOFA-2
COMPONENT fa_inv1impapp
	PORT(b : IN STD_LOGIC;
		 a : IN STD_LOGIC;
		 ci : IN STD_LOGIC;
		 co : OUT STD_LOGIC;
		 s : OUT STD_LOGIC
	);
END COMPONENT;
--Component declaration of AIFA-1
COMPONENT fainvapp
	PORT(b : IN STD_LOGIC;
		 a : IN STD_LOGIC;
		 ci : IN STD_LOGIC;
		 co : OUT STD_LOGIC;
		 s : OUT STD_LOGIC
	);
END COMPONENT;
--Component declaration of EFA
COMPONENT fa_opt2
	PORT(bf : IN STD_LOGIC;
		 af : IN STD_LOGIC;
		 c1 : IN STD_LOGIC;
		 sf : OUT STD_LOGIC;
		 cf : OUT STD_LOGIC
	);
END COMPONENT;
--Component declaration of IIC
COMPONENT fa_inv
	PORT(b : IN STD_LOGIC;
		 a : IN STD_LOGIC;
		 ci : IN STD_LOGIC;
		 co : OUT STD_LOGIC;
		 s : OUT STD_LOGIC
	);
END COMPONENT;
--Component declaration of inverting input half adder
COMPONENT ha_invin1
	PORT(ahc : IN STD_LOGIC;
		 bhc : IN STD_LOGIC;
		 hc : OUT STD_LOGIC;
		 sh : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT ands2
	PORT(i1 : IN STD_LOGIC;
		 i2 : IN STD_LOGIC;
		 o1 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT nots
	PORT(Ai : IN STD_LOGIC;
		 Yi : OUT STD_LOGIC
	);
END COMPONENT;
--Component declaration of half adder
COMPONENT haxor1
	PORT(bh : IN STD_LOGIC;
		 ah : IN STD_LOGIC;
		 hc : OUT STD_LOGIC;
		 sh : OUT STD_LOGIC
	);
END COMPONENT;
--Component declaration of two input xnor
COMPONENT xnorvhdl2
	PORT(i1 : IN STD_LOGIC;
		 i2 : IN STD_LOGIC;
		 o1 : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_79 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_80 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_81 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_82 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_83 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_84 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_85 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_86 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_87 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_88 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_89 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_90 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_91 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_92 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_93 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_95 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_96 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_97 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_98 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_99 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_100 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_101 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_102 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_103 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_104 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_105 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_106 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_107 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_108 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_109 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_110 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_111 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_112 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_113 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_114 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_115 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_116 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_117 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_118 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_119 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_120 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_121 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_122 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_123 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_124 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_125 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_126 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_127 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_128 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_129 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_130 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_131 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_132 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_133 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_134 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_135 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_136 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_137 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_138 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_139 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_140 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_141 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_142 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_143 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_144 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_145 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_146 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_147 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_148 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_149 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_150 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_151 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_152 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_153 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_154 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_155 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_156 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_157 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_158 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_159 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_160 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_161 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_162 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_163 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_164 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_165 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_166 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_167 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_168 :  STD_LOGIC;


BEGIN 



b2v_inst : fa_inv1app
PORT MAP(b => SYNTHESIZED_WIRE_0,
		 a => SYNTHESIZED_WIRE_1,
		 ci => SYNTHESIZED_WIRE_2,
		 s => SYNTHESIZED_WIRE_117,
		 co => SYNTHESIZED_WIRE_50);


b2v_inst1 : fa_inv1app
PORT MAP(b => SYNTHESIZED_WIRE_3,
		 a => SYNTHESIZED_WIRE_4,
		 ci => SYNTHESIZED_WIRE_5,
		 s => SYNTHESIZED_WIRE_48,
		 co => SYNTHESIZED_WIRE_64);


b2v_inst12 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_6,
		 a => SYNTHESIZED_WIRE_7,
		 ci => SYNTHESIZED_WIRE_8,
		 co => SYNTHESIZED_WIRE_97,
		 s => SYNTHESIZED_WIRE_92);


b2v_inst121 : nands2
PORT MAP(i1 => b0,
		 i2 => a6,
		 o1 => SYNTHESIZED_WIRE_29);


b2v_inst125 : nands2
PORT MAP(i1 => b4,
		 i2 => a6,
		 o1 => SYNTHESIZED_WIRE_14);


b2v_inst13 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_9,
		 a => SYNTHESIZED_WIRE_10,
		 ci => SYNTHESIZED_WIRE_11,
		 co => SYNTHESIZED_WIRE_100,
		 s => SYNTHESIZED_WIRE_95);


b2v_inst14 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_12,
		 a => SYNTHESIZED_WIRE_13,
		 ci => SYNTHESIZED_WIRE_14,
		 co => SYNTHESIZED_WIRE_103,
		 s => SYNTHESIZED_WIRE_98);


b2v_inst149 : nands2
PORT MAP(i1 => b1,
		 i2 => a5,
		 o1 => SYNTHESIZED_WIRE_28);


b2v_inst15 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_15,
		 a => SYNTHESIZED_WIRE_16,
		 ci => SYNTHESIZED_WIRE_17,
		 co => SYNTHESIZED_WIRE_123,
		 s => SYNTHESIZED_WIRE_101);


b2v_inst150 : nands2
PORT MAP(i1 => b1,
		 i2 => a6,
		 o1 => SYNTHESIZED_WIRE_46);


b2v_inst151 : nands2
PORT MAP(i1 => b2,
		 i2 => a5,
		 o1 => SYNTHESIZED_WIRE_45);


b2v_inst152 : nands2
PORT MAP(i1 => b2,
		 i2 => a6,
		 o1 => SYNTHESIZED_WIRE_51);


b2v_inst153 : nands2
PORT MAP(i1 => b0,
		 i2 => a5,
		 o1 => SYNTHESIZED_WIRE_21);


b2v_inst154 : nands2
PORT MAP(i1 => b0,
		 i2 => a4,
		 o1 => SYNTHESIZED_WIRE_24);


b2v_inst155 : nands2
PORT MAP(i1 => b0,
		 i2 => a3,
		 o1 => SYNTHESIZED_WIRE_3);


b2v_inst156 : nands2
PORT MAP(i1 => b0,
		 i2 => a2,
		 o1 => SYNTHESIZED_WIRE_0);


b2v_inst157 : nands2
PORT MAP(i1 => b0,
		 i2 => a1,
		 o1 => SYNTHESIZED_WIRE_105);


b2v_inst158 : nands2
PORT MAP(i1 => b1,
		 i2 => a0,
		 o1 => SYNTHESIZED_WIRE_104);


b2v_inst159 : nands2
PORT MAP(i1 => b2,
		 i2 => a0,
		 o1 => SYNTHESIZED_WIRE_2);


b2v_inst160 : nands2
PORT MAP(i1 => b1,
		 i2 => a1,
		 o1 => SYNTHESIZED_WIRE_1);


b2v_inst161 : nands2
PORT MAP(i1 => b1,
		 i2 => a2,
		 o1 => SYNTHESIZED_WIRE_4);


b2v_inst162 : nands2
PORT MAP(i1 => b1,
		 i2 => a3,
		 o1 => SYNTHESIZED_WIRE_25);


b2v_inst163 : nands2
PORT MAP(i1 => b1,
		 i2 => a4,
		 o1 => SYNTHESIZED_WIRE_22);


b2v_inst164 : nands2
PORT MAP(i1 => b2,
		 i2 => a3,
		 o1 => SYNTHESIZED_WIRE_23);


b2v_inst165 : nands2
PORT MAP(i1 => b2,
		 i2 => a4,
		 o1 => SYNTHESIZED_WIRE_27);


b2v_inst166 : nands2
PORT MAP(i1 => b2,
		 i2 => a2,
		 o1 => SYNTHESIZED_WIRE_26);


b2v_inst167 : nands2
PORT MAP(i1 => b2,
		 i2 => a1,
		 o1 => SYNTHESIZED_WIRE_5);


b2v_inst168 : nands2
PORT MAP(i1 => b5,
		 i2 => a5,
		 o1 => SYNTHESIZED_WIRE_13);


b2v_inst169 : nands2
PORT MAP(i1 => b5,
		 i2 => a6,
		 o1 => SYNTHESIZED_WIRE_16);


b2v_inst17 : fainvimpapp
PORT MAP(b => SYNTHESIZED_WIRE_18,
		 a => SYNTHESIZED_WIRE_19,
		 ci => SYNTHESIZED_WIRE_20,
		 co => SYNTHESIZED_WIRE_115,
		 s => SYNTHESIZED_WIRE_163);


b2v_inst170 : nands2
PORT MAP(i1 => b6,
		 i2 => a5,
		 o1 => SYNTHESIZED_WIRE_15);


b2v_inst171 : nands2
PORT MAP(i1 => b6,
		 i2 => a6,
		 o1 => SYNTHESIZED_WIRE_118);


b2v_inst172 : nands2
PORT MAP(i1 => b4,
		 i2 => a5,
		 o1 => SYNTHESIZED_WIRE_11);


b2v_inst173 : nands2
PORT MAP(i1 => b4,
		 i2 => a4,
		 o1 => SYNTHESIZED_WIRE_8);


b2v_inst174 : nands2
PORT MAP(i1 => b4,
		 i2 => a3,
		 o1 => SYNTHESIZED_WIRE_41);


b2v_inst175 : nands2
PORT MAP(i1 => b4,
		 i2 => a2,
		 o1 => SYNTHESIZED_WIRE_32);


b2v_inst176 : nands2
PORT MAP(i1 => b4,
		 i2 => a1,
		 o1 => SYNTHESIZED_WIRE_107);


b2v_inst177 : nands2
PORT MAP(i1 => b5,
		 i2 => a0,
		 o1 => SYNTHESIZED_WIRE_106);


b2v_inst178 : nands2
PORT MAP(i1 => b6,
		 i2 => a0,
		 o1 => SYNTHESIZED_WIRE_30);


b2v_inst179 : nands2
PORT MAP(i1 => b5,
		 i2 => a1,
		 o1 => SYNTHESIZED_WIRE_31);


b2v_inst18 : fa_inv1impapp
PORT MAP(b => SYNTHESIZED_WIRE_21,
		 a => SYNTHESIZED_WIRE_22,
		 ci => SYNTHESIZED_WIRE_23,
		 co => SYNTHESIZED_WIRE_35,
		 s => SYNTHESIZED_WIRE_18);


b2v_inst180 : nands2
PORT MAP(i1 => b5,
		 i2 => a2,
		 o1 => SYNTHESIZED_WIRE_40);


b2v_inst181 : nands2
PORT MAP(i1 => b5,
		 i2 => a3,
		 o1 => SYNTHESIZED_WIRE_7);


b2v_inst182 : nands2
PORT MAP(i1 => b5,
		 i2 => a4,
		 o1 => SYNTHESIZED_WIRE_10);


b2v_inst183 : nands2
PORT MAP(i1 => b6,
		 i2 => a3,
		 o1 => SYNTHESIZED_WIRE_9);


b2v_inst184 : nands2
PORT MAP(i1 => b6,
		 i2 => a4,
		 o1 => SYNTHESIZED_WIRE_12);


b2v_inst185 : nands2
PORT MAP(i1 => b6,
		 i2 => a2,
		 o1 => SYNTHESIZED_WIRE_6);


b2v_inst186 : nands2
PORT MAP(i1 => b6,
		 i2 => a1,
		 o1 => SYNTHESIZED_WIRE_39);


b2v_inst189 : nands2
PORT MAP(i1 => b3,
		 i2 => a0,
		 o1 => SYNTHESIZED_WIRE_49);


b2v_inst190 : nands2
PORT MAP(i1 => b3,
		 i2 => a1,
		 o1 => SYNTHESIZED_WIRE_63);


b2v_inst191 : nands2
PORT MAP(i1 => b3,
		 i2 => a3,
		 o1 => SYNTHESIZED_WIRE_34);


b2v_inst192 : nands2
PORT MAP(i1 => b3,
		 i2 => a2,
		 o1 => SYNTHESIZED_WIRE_19);


b2v_inst194 : nands2
PORT MAP(i1 => b3,
		 i2 => a4,
		 o1 => SYNTHESIZED_WIRE_37);


b2v_inst195 : nands2
PORT MAP(i1 => b3,
		 i2 => a5,
		 o1 => SYNTHESIZED_WIRE_111);


b2v_inst196 : nands2
PORT MAP(i1 => b3,
		 i2 => a6,
		 o1 => SYNTHESIZED_WIRE_86);


b2v_inst197 : nands2
PORT MAP(i1 => b3,
		 i2 => a7,
		 o1 => SYNTHESIZED_WIRE_155);


b2v_inst2 : fa_inv1app
PORT MAP(b => SYNTHESIZED_WIRE_24,
		 a => SYNTHESIZED_WIRE_25,
		 ci => SYNTHESIZED_WIRE_26,
		 s => SYNTHESIZED_WIRE_62,
		 co => SYNTHESIZED_WIRE_20);


b2v_inst20 : fa_inv1impapp
PORT MAP(b => SYNTHESIZED_WIRE_27,
		 a => SYNTHESIZED_WIRE_28,
		 ci => SYNTHESIZED_WIRE_29,
		 co => SYNTHESIZED_WIRE_38,
		 s => SYNTHESIZED_WIRE_33);


b2v_inst21 : fa_inv1impapp
PORT MAP(b => SYNTHESIZED_WIRE_30,
		 a => SYNTHESIZED_WIRE_31,
		 ci => SYNTHESIZED_WIRE_32,
		 co => SYNTHESIZED_WIRE_44,
		 s => SYNTHESIZED_WIRE_125);


b2v_inst22 : fainvimpapp
PORT MAP(b => SYNTHESIZED_WIRE_33,
		 a => SYNTHESIZED_WIRE_34,
		 ci => SYNTHESIZED_WIRE_35,
		 co => SYNTHESIZED_WIRE_132,
		 s => SYNTHESIZED_WIRE_114);


b2v_inst23 : fainvimpapp
PORT MAP(b => SYNTHESIZED_WIRE_36,
		 a => SYNTHESIZED_WIRE_37,
		 ci => SYNTHESIZED_WIRE_38,
		 co => SYNTHESIZED_WIRE_150,
		 s => SYNTHESIZED_WIRE_133);


b2v_inst24 : fa_inv1impapp
PORT MAP(b => SYNTHESIZED_WIRE_39,
		 a => SYNTHESIZED_WIRE_40,
		 ci => SYNTHESIZED_WIRE_41,
		 co => SYNTHESIZED_WIRE_94,
		 s => SYNTHESIZED_WIRE_42);


b2v_inst25 : fainvimpapp
PORT MAP(b => SYNTHESIZED_WIRE_42,
		 a => SYNTHESIZED_WIRE_43,
		 ci => SYNTHESIZED_WIRE_44,
		 co => SYNTHESIZED_WIRE_151,
		 s => SYNTHESIZED_WIRE_142);


b2v_inst26 : fa_inv1impapp
PORT MAP(b => SYNTHESIZED_WIRE_45,
		 a => SYNTHESIZED_WIRE_46,
		 ci => SYNTHESIZED_WIRE_47,
		 co => SYNTHESIZED_WIRE_113,
		 s => SYNTHESIZED_WIRE_36);


b2v_inst3 : fainvapp
PORT MAP(b => SYNTHESIZED_WIRE_48,
		 a => SYNTHESIZED_WIRE_49,
		 ci => SYNTHESIZED_WIRE_50,
		 co => SYNTHESIZED_WIRE_130,
		 s => SYNTHESIZED_WIRE_129);


b2v_inst32 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_51,
		 a => SYNTHESIZED_WIRE_52,
		 ci => Low,
		 co => SYNTHESIZED_WIRE_88,
		 s => SYNTHESIZED_WIRE_112);


b2v_inst37 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_53,
		 af => SYNTHESIZED_WIRE_54,
		 c1 => SYNTHESIZED_WIRE_55,
		 sf => p14,
		 cf => SYNTHESIZED_WIRE_158);


b2v_inst38 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_56,
		 af => SYNTHESIZED_WIRE_57,
		 c1 => SYNTHESIZED_WIRE_58,
		 sf => p13,
		 cf => SYNTHESIZED_WIRE_55);


b2v_inst39 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_59,
		 af => SYNTHESIZED_WIRE_60,
		 c1 => SYNTHESIZED_WIRE_61,
		 sf => p12,
		 cf => SYNTHESIZED_WIRE_58);


b2v_inst4 : fainvapp
PORT MAP(b => SYNTHESIZED_WIRE_62,
		 a => SYNTHESIZED_WIRE_63,
		 ci => SYNTHESIZED_WIRE_64,
		 co => SYNTHESIZED_WIRE_164,
		 s => SYNTHESIZED_WIRE_131);


b2v_inst40 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_65,
		 af => SYNTHESIZED_WIRE_66,
		 c1 => SYNTHESIZED_WIRE_67,
		 sf => p11,
		 cf => SYNTHESIZED_WIRE_61);


b2v_inst41 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_68,
		 af => SYNTHESIZED_WIRE_69,
		 c1 => SYNTHESIZED_WIRE_70,
		 sf => p10,
		 cf => SYNTHESIZED_WIRE_67);


b2v_inst42 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_71,
		 af => SYNTHESIZED_WIRE_72,
		 c1 => SYNTHESIZED_WIRE_73,
		 sf => p9,
		 cf => SYNTHESIZED_WIRE_70);


b2v_inst43 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_74,
		 af => SYNTHESIZED_WIRE_75,
		 c1 => SYNTHESIZED_WIRE_76,
		 sf => p8,
		 cf => SYNTHESIZED_WIRE_73);


b2v_inst44 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_77,
		 af => SYNTHESIZED_WIRE_78,
		 c1 => SYNTHESIZED_WIRE_79,
		 sf => p6,
		 cf => SYNTHESIZED_WIRE_82);


b2v_inst45 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_80,
		 af => SYNTHESIZED_WIRE_81,
		 c1 => SYNTHESIZED_WIRE_82,
		 sf => p7,
		 cf => SYNTHESIZED_WIRE_76);


b2v_inst46 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_83,
		 af => SYNTHESIZED_WIRE_84,
		 c1 => SYNTHESIZED_WIRE_85,
		 sf => SYNTHESIZED_WIRE_65,
		 cf => SYNTHESIZED_WIRE_60);


b2v_inst52 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_86,
		 a => SYNTHESIZED_WIRE_87,
		 ci => SYNTHESIZED_WIRE_88,
		 co => SYNTHESIZED_WIRE_156,
		 s => SYNTHESIZED_WIRE_152);


b2v_inst53 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_89,
		 af => SYNTHESIZED_WIRE_90,
		 c1 => SYNTHESIZED_WIRE_91,
		 sf => SYNTHESIZED_WIRE_68,
		 cf => SYNTHESIZED_WIRE_66);


b2v_inst55 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_92,
		 a => SYNTHESIZED_WIRE_93,
		 ci => SYNTHESIZED_WIRE_94,
		 co => SYNTHESIZED_WIRE_154,
		 s => SYNTHESIZED_WIRE_145);


b2v_inst56 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_95,
		 a => SYNTHESIZED_WIRE_96,
		 ci => SYNTHESIZED_WIRE_97,
		 co => SYNTHESIZED_WIRE_157,
		 s => SYNTHESIZED_WIRE_148);


b2v_inst57 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_98,
		 a => SYNTHESIZED_WIRE_99,
		 ci => SYNTHESIZED_WIRE_100,
		 co => SYNTHESIZED_WIRE_83,
		 s => SYNTHESIZED_WIRE_91);


b2v_inst58 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_101,
		 a => SYNTHESIZED_WIRE_102,
		 ci => SYNTHESIZED_WIRE_103,
		 co => SYNTHESIZED_WIRE_135,
		 s => SYNTHESIZED_WIRE_85);


b2v_inst59 : ha_invin1
PORT MAP(ahc => SYNTHESIZED_WIRE_104,
		 bhc => SYNTHESIZED_WIRE_105,
		 hc => SYNTHESIZED_WIRE_121,
		 sh => p1);


b2v_inst60 : ha_invin1
PORT MAP(ahc => SYNTHESIZED_WIRE_106,
		 bhc => SYNTHESIZED_WIRE_107,
		 hc => SYNTHESIZED_WIRE_126,
		 sh => SYNTHESIZED_WIRE_160);


b2v_inst61 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_108,
		 a => SYNTHESIZED_WIRE_109,
		 ci => SYNTHESIZED_WIRE_110,
		 co => SYNTHESIZED_WIRE_139,
		 s => SYNTHESIZED_WIRE_136);


b2v_inst62 : ands2
PORT MAP(i1 => b7,
		 i2 => a7,
		 o1 => SYNTHESIZED_WIRE_138);


b2v_inst63 : ands2
PORT MAP(i1 => b0,
		 i2 => a7,
		 o1 => SYNTHESIZED_WIRE_47);


b2v_inst64 : ands2
PORT MAP(i1 => b1,
		 i2 => a7,
		 o1 => SYNTHESIZED_WIRE_52);


b2v_inst65 : ands2
PORT MAP(i1 => b2,
		 i2 => a7,
		 o1 => SYNTHESIZED_WIRE_87);


b2v_inst66 : ands2
PORT MAP(i1 => b4,
		 i2 => a7,
		 o1 => SYNTHESIZED_WIRE_17);


b2v_inst67 : ands2
PORT MAP(i1 => b5,
		 i2 => a7,
		 o1 => SYNTHESIZED_WIRE_119);


b2v_inst68 : ands2
PORT MAP(i1 => b6,
		 i2 => a7,
		 o1 => SYNTHESIZED_WIRE_109);


b2v_inst69 : fa_inv
PORT MAP(b => SYNTHESIZED_WIRE_111,
		 a => SYNTHESIZED_WIRE_112,
		 ci => SYNTHESIZED_WIRE_113,
		 co => SYNTHESIZED_WIRE_153,
		 s => SYNTHESIZED_WIRE_149);


b2v_inst7 : ands2
PORT MAP(i1 => b0,
		 i2 => a0,
		 o1 => p0);


b2v_inst70 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_114,
		 af => SYNTHESIZED_WIRE_115,
		 c1 => SYNTHESIZED_WIRE_116,
		 sf => SYNTHESIZED_WIRE_77,
		 cf => SYNTHESIZED_WIRE_81);


b2v_inst71 : nots
PORT MAP(Ai => SYNTHESIZED_WIRE_117,
		 Yi => SYNTHESIZED_WIRE_122);


b2v_inst72 : fa_inv1
PORT MAP(b => SYNTHESIZED_WIRE_118,
		 a => SYNTHESIZED_WIRE_119,
		 ci => SYNTHESIZED_WIRE_120,
		 co => SYNTHESIZED_WIRE_110,
		 s => SYNTHESIZED_WIRE_124);


b2v_inst73 : haxor1
PORT MAP(bh => SYNTHESIZED_WIRE_121,
		 ah => SYNTHESIZED_WIRE_122,
		 hc => SYNTHESIZED_WIRE_128,
		 sh => p2);


b2v_inst74 : ha_invin1
PORT MAP(ahc => SYNTHESIZED_WIRE_123,
		 bhc => SYNTHESIZED_WIRE_124,
		 hc => SYNTHESIZED_WIRE_137,
		 sh => SYNTHESIZED_WIRE_134);


b2v_inst75 : nots
PORT MAP(Ai => SYNTHESIZED_WIRE_125,
		 Yi => SYNTHESIZED_WIRE_127);


b2v_inst76 : haxor1
PORT MAP(bh => SYNTHESIZED_WIRE_126,
		 ah => SYNTHESIZED_WIRE_127,
		 hc => SYNTHESIZED_WIRE_141,
		 sh => SYNTHESIZED_WIRE_78);


b2v_inst77 : haxor1
PORT MAP(bh => SYNTHESIZED_WIRE_128,
		 ah => SYNTHESIZED_WIRE_129,
		 hc => SYNTHESIZED_WIRE_168,
		 sh => p3);


b2v_inst78 : haxor1
PORT MAP(bh => SYNTHESIZED_WIRE_130,
		 ah => SYNTHESIZED_WIRE_131,
		 hc => SYNTHESIZED_WIRE_165,
		 sh => SYNTHESIZED_WIRE_166);


b2v_inst79 : haxor1
PORT MAP(bh => SYNTHESIZED_WIRE_132,
		 ah => SYNTHESIZED_WIRE_133,
		 hc => SYNTHESIZED_WIRE_144,
		 sh => SYNTHESIZED_WIRE_140);


b2v_inst8 : ands2
PORT MAP(i1 => b4,
		 i2 => a0,
		 o1 => SYNTHESIZED_WIRE_167);


b2v_inst80 : haxor1
PORT MAP(bh => SYNTHESIZED_WIRE_134,
		 ah => SYNTHESIZED_WIRE_135,
		 hc => SYNTHESIZED_WIRE_57,
		 sh => SYNTHESIZED_WIRE_59);


b2v_inst81 : haxor1
PORT MAP(bh => SYNTHESIZED_WIRE_136,
		 ah => SYNTHESIZED_WIRE_137,
		 hc => SYNTHESIZED_WIRE_54,
		 sh => SYNTHESIZED_WIRE_56);


b2v_inst82 : haxor1
PORT MAP(bh => SYNTHESIZED_WIRE_138,
		 ah => SYNTHESIZED_WIRE_139,
		 hc => SYNTHESIZED_WIRE_159,
		 sh => SYNTHESIZED_WIRE_53);


b2v_inst83 : ands2
PORT MAP(i1 => b7,
		 i2 => a6,
		 o1 => SYNTHESIZED_WIRE_108);


b2v_inst84 : ands2
PORT MAP(i1 => b7,
		 i2 => a5,
		 o1 => SYNTHESIZED_WIRE_120);


b2v_inst85 : ands2
PORT MAP(i1 => b7,
		 i2 => a4,
		 o1 => SYNTHESIZED_WIRE_102);


b2v_inst86 : ands2
PORT MAP(i1 => b7,
		 i2 => a3,
		 o1 => SYNTHESIZED_WIRE_99);


b2v_inst87 : ands2
PORT MAP(i1 => b7,
		 i2 => a2,
		 o1 => SYNTHESIZED_WIRE_96);


b2v_inst88 : ands2
PORT MAP(i1 => b7,
		 i2 => a1,
		 o1 => SYNTHESIZED_WIRE_93);


b2v_inst89 : ands2
PORT MAP(i1 => b7,
		 i2 => a0,
		 o1 => SYNTHESIZED_WIRE_43);


b2v_inst90 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_140,
		 af => SYNTHESIZED_WIRE_141,
		 c1 => SYNTHESIZED_WIRE_142,
		 sf => SYNTHESIZED_WIRE_80,
		 cf => SYNTHESIZED_WIRE_75);


b2v_inst91 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_143,
		 af => SYNTHESIZED_WIRE_144,
		 c1 => SYNTHESIZED_WIRE_145,
		 sf => SYNTHESIZED_WIRE_74,
		 cf => SYNTHESIZED_WIRE_72);


b2v_inst92 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_146,
		 af => SYNTHESIZED_WIRE_147,
		 c1 => SYNTHESIZED_WIRE_148,
		 sf => SYNTHESIZED_WIRE_71,
		 cf => SYNTHESIZED_WIRE_69);


b2v_inst93 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_149,
		 af => SYNTHESIZED_WIRE_150,
		 c1 => SYNTHESIZED_WIRE_151,
		 sf => SYNTHESIZED_WIRE_143,
		 cf => SYNTHESIZED_WIRE_147);


b2v_inst94 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_152,
		 af => SYNTHESIZED_WIRE_153,
		 c1 => SYNTHESIZED_WIRE_154,
		 sf => SYNTHESIZED_WIRE_146,
		 cf => SYNTHESIZED_WIRE_90);


b2v_inst95 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_155,
		 af => SYNTHESIZED_WIRE_156,
		 c1 => SYNTHESIZED_WIRE_157,
		 sf => SYNTHESIZED_WIRE_89,
		 cf => SYNTHESIZED_WIRE_84);


b2v_inst96 : xnorvhdl2
PORT MAP(i1 => SYNTHESIZED_WIRE_158,
		 i2 => SYNTHESIZED_WIRE_159,
		 o1 => p15);


b2v_inst97 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_160,
		 af => SYNTHESIZED_WIRE_161,
		 c1 => SYNTHESIZED_WIRE_162,
		 sf => p5,
		 cf => SYNTHESIZED_WIRE_79);


b2v_inst98 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_163,
		 af => SYNTHESIZED_WIRE_164,
		 c1 => SYNTHESIZED_WIRE_165,
		 sf => SYNTHESIZED_WIRE_161,
		 cf => SYNTHESIZED_WIRE_116);


b2v_inst99 : fa_opt2
PORT MAP(bf => SYNTHESIZED_WIRE_166,
		 af => SYNTHESIZED_WIRE_167,
		 c1 => SYNTHESIZED_WIRE_168,
		 sf => p4,
		 cf => SYNTHESIZED_WIRE_162);


END bdf_type;
